module instruction_mem #(
    parameter MEM_SIZE = 58
)
(
   input  logic [31:0] addr,
   output logic [31:0] data
);

   // Read-memory that contains all RV32I instructions
   logic [31:0] instrs [MEM_SIZE];
   assign instrs = {{12'b10101, 5'd0, 3'b000, 5'd1, 7'b0010011}, 
                    {12'b111, 5'd0, 3'b000, 5'd2, 7'b0010011}, 
                    {12'b111111111100, 5'd0, 3'b000, 5'd3, 7'b0010011}, 
                    {12'b1011100, 5'd1, 3'b111, 5'd5, 7'b0010011}, 
                    {12'b10101, 5'd5, 3'b100, 5'd5, 7'b0010011}, 
                    {12'b1011100, 5'd1, 3'b110, 5'd6, 7'b0010011}, 
                    {12'b1011100, 5'd6, 3'b100, 5'd6, 7'b0010011}, 
                    {12'b111, 5'd1, 3'b000, 5'd7, 7'b0010011}, 
                    {12'b11101, 5'd7, 3'b100, 5'd7, 7'b0010011}, 
                    {6'b000000, 6'b110, 5'd1, 3'b001, 5'd8, 7'b0010011}, 
                    {12'b10101000001, 5'd8, 3'b100, 5'd8, 7'b0010011}, 
                    {6'b000000, 6'b10, 5'd1, 3'b101, 5'd9, 7'b0010011}, 
                    {12'b100, 5'd9, 3'b100, 5'd9, 7'b0010011}, 
                    {7'b0000000, 5'd2, 5'd1, 3'b111, 5'd10, 7'b0110011}, 
                    {12'b100, 5'd10, 3'b100, 5'd10, 7'b0010011}, 
                    {7'b0000000, 5'd2, 5'd1, 3'b110, 5'd11, 7'b0110011}, 
                    {12'b10110, 5'd11, 3'b100, 5'd11, 7'b0010011}, 
                    {7'b0000000, 5'd2, 5'd1, 3'b100, 5'd12, 7'b0110011}, 
                    {12'b10011, 5'd12, 3'b100, 5'd12, 7'b0010011}, 
                    {7'b0000000, 5'd2, 5'd1, 3'b000, 5'd13, 7'b0110011}, 
                    {12'b11101, 5'd13, 3'b100, 5'd13, 7'b0010011}, 
                    {7'b0100000, 5'd2, 5'd1, 3'b000, 5'd14, 7'b0110011}, 
                    {12'b1111, 5'd14, 3'b100, 5'd14, 7'b0010011}, 
                    {7'b0000000, 5'd2, 5'd2, 3'b001, 5'd15, 7'b0110011}, 
                    {12'b1110000001, 5'd15, 3'b100, 5'd15, 7'b0010011}, 
                    {7'b0000000, 5'd2, 5'd1, 3'b101, 5'd16, 7'b0110011}, 
                    {12'b1, 5'd16, 3'b100, 5'd16, 7'b0010011}, 
                    {7'b0000000, 5'd1, 5'd2, 3'b011, 5'd17, 7'b0110011}, 
                    {12'b0, 5'd17, 3'b100, 5'd17, 7'b0010011}, 
                    {12'b10101, 5'd2, 3'b011, 5'd18, 7'b0010011}, 
                    {12'b0, 5'd18, 3'b100, 5'd18, 7'b0010011}, 
                    {20'b00000000000000000000, 5'd19, 7'b0110111}, 
                    {12'b1, 5'd19, 3'b100, 5'd19, 7'b0010011}, 
                    {6'b010000, 6'b1, 5'd3, 3'b101, 5'd20, 7'b0010011}, 
                    {12'b111111111111, 5'd20, 3'b100, 5'd20, 7'b0010011}, 
                    {7'b0000000, 5'd1, 5'd3, 3'b010, 5'd21, 7'b0110011}, 
                    {12'b0, 5'd21, 3'b100, 5'd21, 7'b0010011}, 
                    {12'b1, 5'd3, 3'b010, 5'd22, 7'b0010011}, 
                    {12'b0, 5'd22, 3'b100, 5'd22, 7'b0010011}, 
                    {7'b0100000, 5'd2, 5'd1, 3'b101, 5'd23, 7'b0110011}, 
                    {12'b1, 5'd23, 3'b100, 5'd23, 7'b0010011}, 
                    {20'b00000000000000000100, 5'd4, 7'b0010111}, 
                    {6'b000000, 6'b111, 5'd4, 3'b101, 5'd24, 7'b0010011}, 
                    {12'b10000000, 5'd24, 3'b100, 5'd24, 7'b0010011}, 
                    {1'b0, 10'b0000000010, 1'b0, 8'b00000000, 5'd25, 7'b1101111}, 
                    {20'b00000000000000000000, 5'd4, 7'b0010111}, 
                    {7'b0000000, 5'd4, 5'd25, 3'b100, 5'd25, 7'b0110011}, 
                    {12'b1, 5'd25, 3'b100, 5'd25, 7'b0010011}, 
                    {12'b10000, 5'd4, 3'b000, 5'd26, 7'b1100111}, 
                    {7'b0100000, 5'd4, 5'd26, 3'b000, 5'd26, 7'b0110011}, 
                    {12'b111111110001, 5'd26, 3'b000, 5'd26, 7'b0010011}, 
                    {7'b0000000, 5'd1, 5'd2, 3'b010, 5'b00001, 7'b0100011}, 
                    {12'b1, 5'd2, 3'b010, 5'd27, 7'b0000011}, 
                    {12'b10100, 5'd27, 3'b100, 5'd27, 7'b0010011}, 
                    {12'b1, 5'd0, 3'b000, 5'd28, 7'b0010011}, 
                    {12'b1, 5'd0, 3'b000, 5'd29, 7'b0010011}, 
                    {12'b1, 5'd0, 3'b000, 5'd30, 7'b0010011}, 
                    {1'b0, 10'b0000000000, 1'b0, 8'b00000000, 5'd0, 7'b1101111}};
	assign data = instrs[addr[$clog2($size(instrs)) + 1 : 2]];
	
endmodule
