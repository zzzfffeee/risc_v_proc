/* RISC-V CPU Core defines */
`define DATA_WIDTH 32
`define DATA_MEM_SIZE 32
`define PROG_MEM_SIZE 58
`define NUM_CORE_REGS 31
